`timescale 1ns/10ps

module control_unit_tb;




endmodule

